module alu(
  input wire [31:0] op1, // rs1;
  input wire [31:0] op2, // rs2 or Immediate;
  input wire [31:0] instr, // instruction
  output reg [31:0] res); // result 




endmodule